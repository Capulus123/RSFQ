
.subckt THmitll_AND2 a b clk q
.model jjmit jj(rtype=1, vg=2.8mV, cap=0.07pF, r0=160, rn=16, icrit=0.1mA)
.param Phi0=2.067833848E-15
.param B0=1
.param Ic0=0.0001
.param IcRs=100u*6.859904418
.param B0Rs=IcRs/Ic0*B0
.param Rsheet=2 
.param Lsheet=1.13e-12 
.param LP=0.5p
.param IC=2.5
.param LB=2p
.param BiasCoef=0.7
.param B1=2.5
.param B2=1.60
.param B3=1.94
.param B4=1.57
.param B5=1.25
.param B6=1.25
.param B7=2.5
.param B8=1.60
.param B9=1.94
.param B10=1.57
.param B11=1.25
.param B12=1.25
.param B13=2.5
.param B14=1.71
.param B15=2.5
.param IB1=175u
.param IB2=162u
.param IB3=175u
.param IB4=162u
.param IB5=175u
.param IB6=124u
.param IB7=175u
.param LB1=LB
.param LB2=LB
.param LB3=LB
.param LB4=LB
.param LB5=LB
.param LB6=LB
.param LB7=LB
.param L1=1.8843p
.param L2=4.2266p
.param L3=9.6820p
.param L4=0.9913p
.param L5=2.5745p
.param L6=1.8843p
.param L7=4.2266p
.param L8=9.6820p
.param L9=0.9913p
.param L10=2.5745p
.param L11=1.5293p
.param L12=2.6230p
.param L13=0.7965p
.param L14=0.7671p
.param L15=1.2144p
.param LP1=LP
.param LP3=LP
.param LP4=LP
.param LP7=LP
.param LP9=LP
.param LP10=LP
.param LP13=LP
.param LP14=LP
.param LP15=LP
.param RB1=B0Rs/B1
.param RB2=B0Rs/B2
.param RB3=B0Rs/B3
.param RB4=B0Rs/B4
.param RB5=B0Rs/B5
.param RB6=B0Rs/B6
.param RB7=B0Rs/B7
.param RB8=B0Rs/B8
.param RB9=B0Rs/B9
.param RB10=B0Rs/B10
.param RB11=B0Rs/B11
.param RB12=B0Rs/B12
.param RB13=B0Rs/B13
.param RB14=B0Rs/B14
.param RB15=B0Rs/B15
.param LRB1=(RB1/Rsheet)*Lsheet+LP
.param LRB2=(RB2/Rsheet)*Lsheet
.param LRB3=(RB3/Rsheet)*Lsheet+LP
.param LRB4=(RB4/Rsheet)*Lsheet+LP
.param LRB5=(RB5/Rsheet)*Lsheet
.param LRB6=(RB6/Rsheet)*Lsheet
.param LRB7=(RB7/Rsheet)*Lsheet+LP
.param LRB8=(RB8/Rsheet)*Lsheet
.param LRB9=(RB9/Rsheet)*Lsheet+LP
.param LRB10=(RB10/Rsheet)*Lsheet+LP
.param LRB11=(RB11/Rsheet)*Lsheet
.param LRB12=(RB12/Rsheet)*Lsheet
.param LRB13=(RB13/Rsheet)*Lsheet+LP
.param LRB14=(RB14/Rsheet)*Lsheet+LP
.param LRB15=(RB15/Rsheet)*Lsheet+LP
B1 1 2 jjmit  area=B1 
B2 4 5 jjmit  area=B2 
B3 5 6 jjmit  area=B3 
B4 8 9 jjmit  area=B4 
B5 8 10 jjmit  area=B5 
B6 12 13 jjmit  area=B6 
B7 14 15 jjmit  area=B7 
B8 17 18 jjmit  area=B8 
B9 18 19 jjmit  area=B9 
B10 21 22 jjmit  area=B10 
B11 21 23 jjmit  area=B11 
B12 24 13 jjmit  area=B12 
B13 25 26 jjmit  area=B13 
B14 28 29 jjmit  area=B14 
B15 31 32 jjmit  area=B15
IB1 0 3 pwl(0 0 5p IB1)
IB2 0 7 pwl(0 0 5p IB2)
IB3 0 16 pwl(0 0 5p IB3)
IB4 0 20 pwl(0 0 5p IB4)
IB5 0 27 pwl(0 0 5p IB5)
IB6 0 30 pwl(0 0 5p IB6)
IB7 0 33 pwl(0 0 5p IB7)
LB1 3 1 1.032E-012 
LB2 7 5 3.135E-012 
LB3 16 14 1.016E-012 
LB4 20 18 3.19E-012 
LB5 27 25 1.708E-012 
LB6 30 28 6.363E-013 
LB7 33 31 7.55E-013 
L1 a 1 1.874E-012 
L2 1 4 4.249E-012 
L3 5 8 9.672E-012 
L4 10 11 9.976E-013 
L5 8 12 2.561E-012 
L6 b 14 1.875E-012 
L7 14 17 4.233E-012 
L8 18 21 9.691E-012 
L9 11 23 9.928E-013 
L10 21 24 2.556E-012 
L11 clk 25 1.531E-012 
L12 25 28 2.626E-012 
L13 28 11 7.973E-013 
L14 13 31 7.691E-013 
L15 31 q 1.217E-012 
LP1 2 0 3.464E-013 
LP3 6 0 6.827E-013 
LP4 0 9 4.723E-013 
LP7 15 0 3.484E-013 
LP9 19 0 6.81E-013 
LP10 22 0 4.756E-013 
LP13 26 0 3.392E-013 
LP14 29 0 3.972E-013 
LP15 32 0 3.699E-013 
RB1 1 101 RB1  
LRB1 101 0 LRB1 
RB2 4 104 RB2  
LRB2 104 5 LRB2 
RB3 5 105 RB3  
LRB3 105 0 LRB3 
RB4 108 8 RB4  
LRB4 0 108 LRB4 
RB5 8 110 RB5  
LRB5 110 10 LRB5 
RB6 12 112 RB6  
LRB6 112 13 LRB6 
RB7 14 114 RB7  
LRB7 114 0 LRB7 
RB8 17 117 RB8  
LRB8 117 18 LRB8 
RB9 18 118 RB9  
LRB9 118 0 LRB9 
RB10 21 121 RB10  
LRB10 121 0 LRB10 
RB11 123 21 RB11  
LRB11 23 123 LRB11 
RB12 24 124 RB12  
LRB12 124 13 LRB12 
RB13 25 125 RB13  
LRB13 125 0 LRB13 
RB14 28 128 RB14  
LRB14 128 0 LRB14 
RB15 31 131 RB15  
LRB15 131 0 LRB15 
.ends

* === SOURCE DEFINITION ===

.subckt SOURCECELL  a q
.model jjmit jj(rtype=1, vg=2.8mv, cap=0.07pf, r0=160, rn=16, icrit=0.1ma)
.param phi0=2.067833848e-15
.param b0=1
.param ic0=0.0001
.param icrs=100u*6.859904418
.param b0rs=icrs/ic0*b0
.param rsheet=2
.param lsheet=1.13e-12
.param lp=0.5p
.param ic=2.5
.param lb=2p
.param biascoef=0.7
.param b1=2.25
.param b2=2.25
.param b3=ic
.param ib1=275u
.param ib2=b3*ic0*biascoef
.param lb1=lb
.param lb2=lb
.param l1=1p
.param l2=3.9p
.param l3=0.6p
.param l4=1.1p
.param l5=4.5p
.param l6=phi0/(4*ic*ic0)
.param lp2=lp
.param lp3=lp
.param rb1=b0rs/b1
.param rb2=b0rs/b2
.param rb3=b0rs/b3
.param lrb1=(rb1/rsheet)*lsheet
.param lrb2=(rb2/rsheet)*lsheet+lp
.param lrb3=(rb3/rsheet)*lsheet+lp
b1 2 3 jjmit  area=b1
b2 5 6 jjmit  area=b2
b3 7 8 jjmit  area=b3
ib1 0 4 pwl(0 0 5p ib1)
ib2 0 9 pwl(0 0 5p ib2)
lb1 4 3 2.825e-012
lb2 9 7 2.942e-012
l1 a 1 1.672e-012
l2 1 0 3.901e-012
l3 1 2 5.953e-013
l4 3 5 1.1e-012
l5 5 7 4.542e-012
l6 7 q 2.012e-012
lp2 6 0 3.924e-013
lp3 8 0 3.841e-013
rb1 2 102 rb1
lrb1 102 3 lrb1
rb2 5 105 rb2
lrb2 105 0 lrb2
rb3 7 107 rb3
lrb3 107 0 lrb3
.ends SOURCECELL

* === INPUT LOAD DEFINITION ===

.subckt LOADINCELL  a q
.model jjmit jj(rtype=1, vg=2.8mv, cap=0.07pf, r0=160, rn=16, icrit=0.1ma)
.param phi0=2.067833848e-15
.param b0=1
.param ic0=0.0001
.param icrs=100u*6.859904418
.param b0rs=icrs/ic0*b0
.param rsheet=2
.param lsheet=1.13e-12
.param lp=0.5p
.param ic=2.5
.param lb=2p
.param biascoef=0.7
.param b1=ic
.param b2=ic
.param ib1=(b1+b2)*ic0*biascoef
.param lb1=lb
.param l1=phi0/(4*b1*ic0)
.param l2=phi0/(4*b1*ic0)
.param l3=phi0/(4*b2*ic0)
.param l4=phi0/(4*b2*ic0)
.param lp1=lp
.param lp2=lp
.param rb1=b0rs/b1
.param rb2=b0rs/b2
.param lrb1=(rb1/rsheet)*lsheet+lp
.param lrb2=(rb2/rsheet)*lsheet+lp
b1 1 2 jjmit  area=b1
b2 5 6 jjmit  area=b2
ib1 0 4 pwl(0 0 5p ib1)
lb1 4 3 2.336e-012
l1 a 1 2.07e-012
l2 1 3 2.088e-012
l3 3 5 2.082e-012
l4 5 q 2.072e-012
lp1 2 0 3.137e-013
lp2 6 0 3.123e-013
rb1 1 101 rb1
lrb1 101 0 lrb1
rb2 5 105 rb2
lrb2 105 0 lrb2
.ends LOADINCELL

* === OUTPUT LOAD DEFINITION ===

.subckt LOADOUTCELL  a q
.model jjmit jj(rtype=1, vg=2.8mv, cap=0.07pf, r0=160, rn=16, icrit=0.1ma)
.param phi0=2.067833848e-15
.param b0=1
.param ic0=0.0001
.param icrs=100u*6.859904418
.param b0rs=icrs/ic0*b0
.param rsheet=2
.param lsheet=1.13e-12
.param lp=0.5p
.param ic=2.5
.param lb=2p
.param biascoef=0.7
.param b1=ic
.param b2=ic
.param ib1=(b1+b2)*ic0*biascoef
.param lb1=lb
.param l1=phi0/(4*b1*ic0)
.param l2=phi0/(4*b1*ic0)
.param l3=phi0/(4*b2*ic0)
.param l4=phi0/(4*b2*ic0)
.param lp1=lp
.param lp2=lp
.param rb1=b0rs/b1
.param rb2=b0rs/b2
.param lrb1=(rb1/rsheet)*lsheet+lp
.param lrb2=(rb2/rsheet)*lsheet+lp
b1 1 2 jjmit  area=b1
b2 5 6 jjmit  area=b2
ib1 0 4 pwl(0 0 5p ib1)
lb1 4 3 2.336e-012
l1 a 1 2.07e-012
l2 1 3 2.088e-012
l3 3 5 2.082e-012
l4 5 q 2.072e-012
lp1 2 0 3.137e-013
lp2 6 0 3.123e-013
rb1 1 101 rb1
lrb1 101 0 lrb1
rb2 5 105 rb2
lrb2 105 0 lrb2
.ends LOADOUTCELL

* === SINK DEFINITION ===

.subckt SINKCELL  1
r1 1 0 2
.ends SINKCELL

* ===== MAIN =====

I_a 0 1 pwl(0 0 150p 0 153p 600u 156p 0 250p 0 253p 600u 256p 0 280p 0 283p 600u 286p 0 540p 0 543p 600u 546p 0 600p 0 603p 600u 606p 0 640p 0 643p 600u 646p 0 780p 0 783p 600u 786p 0)
XSOURCEINa 1 2 SOURCECELL
XLOADINa 2 3 LOADINCELL
I_b 0 4 pwl(0 0 350p 0 353p 600u 356p 0 450p 0 453p 600u 456p 0 480p 0 483p 600u 486p 0 560p 0 563p 600u 566p 0 580p 0 583p 600u 586p 0 660p 0 663p 600u 666p 0 740p 0 743p 600u 746p 0)
XSOURCEINb 4 5 SOURCECELL
XLOADINb 5 6 LOADINCELL
I_clk 0 7 pulse(0 600u 20p 2p 2p 1p 100p)
XSOURCEINclk 7 8 SOURCECELL
XLOADINclk 8 9 LOADINCELL
XLOADOUTq 10 11 LOADOUTCELL
XSINKOUTq 11 SINKCELL
XDUT 3 6 9 10 THmitll_AND2
.tran 1p 1000p
.end
